** Profile: "SCHEMATIC1-MC"  [ e:\fuckultate\an ii\sem ii\biggest shit in the world\proiect pwm\version_3\varianta_3-PSpiceFiles\SCHEMATIC1\MC.sim ] 

** Creating circuit file "MC.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\Teo\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 800us 0 100us 
.MC 5 TRAN V([OUT]) YMAX OUTPUT ALL SEED=200 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
