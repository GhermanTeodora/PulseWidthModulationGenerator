** Profile: "SCHEMATIC1-trial2"  [ e:\fuckultate\an ii\sem ii\biggest shit in the world\proiect pwm\version_3\varianta_3-PSpiceFiles\SCHEMATIC1\trial2.sim ] 

** Creating circuit file "trial2.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\Teo\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 800us 0 
.STEP LIN PARAM set20 0 1 0.25 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
